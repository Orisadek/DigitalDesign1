//
// Verilog Module Ori_Alon_Lab_1_lib.control_module
//
// Created:
//          by - orisad.UNKNOWN (TOMER)
//          at - 19:20:41 01/21/2024
//
// using Mentor Graphics HDL Designer(TM) 2019.2 (Build 5)
//

`resetall
`timescale 1ns/10ps
module control_module;


// ### Please start your Verilog code here ### 

endmodule
